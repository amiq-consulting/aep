/******************************************************************************
Copyright (c) 2004-2017, AMIQ Consulting srl. All rights reserved.

Licensed under the Apache License, Version 2.0 (the "License");
you may not use this file except in compliance with the License.
You may obtain a copy of the License at
    http://www.apache.org/licenses/LICENSE-2.0

Unless required by applicable law or agreed to in writing, software
distributed under the License is distributed on an "AS IS" BASIS,
WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
See the License for the specific language governing permissions and
limitations under the License.
 *******************************************************************************/
 
`ifndef __ex_out_monitor
`define __ex_out_monitor

/**
 * TODO: declare the ex_out_monitor class 
 * 
 * 
 * TODO: declare a virtual interface ex_out_intf field
 * 
 * 
 * TODO: declare a field of type ex_out_serial_obj
 * 
 * 
 * TODO: declare an event new_cmd_e
 * 
 * TODO: implement a task monitor() that recovers the data transfers from the serial bus and translates them into ex_out_serial_obj
 * This task should be sensitive to reset and wait for the release of reset before starting collecting items on the bus.
 * 
 * 
 */

`endif


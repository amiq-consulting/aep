
/******************************************************************************
Copyright (c) 2004-2017, AMIQ Consulting srl. All rights reserved.

Licensed under the Apache License, Version 2.0 (the "License");
you may not use this file except in compliance with the License.
You may obtain a copy of the License at
    http://www.apache.org/licenses/LICENSE-2.0

Unless required by applicable law or agreed to in writing, software
distributed under the License is distributed on an "AS IS" BASIS,
WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
See the License for the specific language governing permissions and
limitations under the License.
 *******************************************************************************/

`ifndef __ex_out_pkg
`define __ex_out_pkg

/**
 * TODO: declare package ex_pkg
 * 
 * 
 * TODO: import ex_in_pkg and ex_out_pkg
 * 
 * 
 * TODO: inside ex_pkg include all ex_* files
**/


`endif




/******************************************************************************
Copyright (c) 2004-2017, AMIQ Consulting srl. All rights reserved.

Licensed under the Apache License, Version 2.0 (the "License");
you may not use this file except in compliance with the License.
You may obtain a copy of the License at
    http://www.apache.org/licenses/LICENSE-2.0

Unless required by applicable law or agreed to in writing, software
distributed under the License is distributed on an "AS IS" BASIS,
WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
See the License for the specific language governing permissions and
limitations under the License.
 *******************************************************************************/

`ifndef __ex_in_driver
`define __ex_in_driver

/***
 * TODO: declare the driver class ex_in_driver
 * 
 * 
 * TODO: declare a virtual interface ex_in_intf field inside the driver class 
 * 
 * 
 * TODO: declare a task drive_command(ex_in_cmd acmd) which drives the argument on input wires
 * 
 * 
 * TODO: declare a task scenario() that creates 10 commands and drives them on the bus using the drive_command() task
 * This task should be sensitive to reset and wait for the release of reset before starting to drive items.
 * 
 * 
 * 
**/

`endif

/******************************************************************************
Copyright (c) 2004-2017, AMIQ Consulting srl. All rights reserved.

Licensed under the Apache License, Version 2.0 (the "License");
you may not use this file except in compliance with the License.
You may obtain a copy of the License at
    http://www.apache.org/licenses/LICENSE-2.0

Unless required by applicable law or agreed to in writing, software
distributed under the License is distributed on an "AS IS" BASIS,
WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
See the License for the specific language governing permissions and
limitations under the License.
 *******************************************************************************/
 
`ifndef __ex_in_intf
`define __ex_in_intf

/**
 * 
 * TODO: create the input interface ex_input_intf containing the following port
 * input clk     - 1 bit
 * input reset   - 1 bit
 * 
 * 
 * TODO: declare the following fields inside the input interface
 * addr    - 8 bit
 * data_in - 8 bit
 * rnw     - 1 bit
 * cmd     - 1 bit
 * busy    - 1 bit
**/

`endif
 

/******************************************************************************
Copyright (c) 2004-2017, AMIQ Consulting srl. All rights reserved.

Licensed under the Apache License, Version 2.0 (the "License");
you may not use this file except in compliance with the License.
You may obtain a copy of the License at
    http://www.apache.org/licenses/LICENSE-2.0

Unless required by applicable law or agreed to in writing, software
distributed under the License is distributed on an "AS IS" BASIS,
WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
See the License for the specific language governing permissions and
limitations under the License.
 *******************************************************************************/

`ifndef __ex_in_monitor
`define __ex_in_monitor

/***
 * TODO: declare the monitor class ex_in_monitor
 * 
 * 
 * TODO: declare a virtual interface ex_in_intf field inside the monitor class 
 * 
 * 
 * TODO: declare a field of type ex_in_cmd 
 * 
 * TODO: declare an event new_cmd_e
 * 
 * TODO: declare a task monitor_bus() which recovers data from the wires.
 * This task should be sensitive to reset and wait for the release of reset before starting collecting commands on the bus. 
 * The recovered data is saved into the previously defined field and new data is announced using new_cmd_e 
 *  
 * TODO: declare a functional coverage group that samples the recovered commands parameters
 * 
**/

`endif

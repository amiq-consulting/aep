/******************************************************************************
 Copyright (c) 2004-2018, AMIQ Consulting srl. All rights reserved.

 Licensed under the Apache License, Version 2.0 (the "License");
 you may not use this file except in compliance with the License.
 You may obtain a copy of the License at
 http://www.apache.org/licenses/LICENSE-2.0

 Unless required by applicable law or agreed to in writing, software
 distributed under the License is distributed on an "AS IS" BASIS,
 WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 See the License for the specific language governing permissions and
 limitations under the License.
 *******************************************************************************/

`ifndef __EX_TEST_PKG
`define __EX_TEST_PKG

package ex_test_pkg;


	`include "uvm_macros.svh"
	import uvm_pkg::*;

	import ex_in_pkg::*;
	import ex_out_pkg::*;
	import ex_pkg::*;

	`include "ex_test.svh"


endpackage : ex_test_pkg




`endif


/******************************************************************************
Copyright (c) 2004-2017, AMIQ Consulting srl. All rights reserved.

Licensed under the Apache License, Version 2.0 (the "License");
you may not use this file except in compliance with the License.
You may obtain a copy of the License at
    http://www.apache.org/licenses/LICENSE-2.0

Unless required by applicable law or agreed to in writing, software
distributed under the License is distributed on an "AS IS" BASIS,
WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
See the License for the specific language governing permissions and
limitations under the License.
 *******************************************************************************/

`timescale 1ns/1ns

// TODO: include source files

module ex_top();
   
 // TODO: declare reset, clock and interface specific signals
  
 // TODO: implement a clock generator
 // TODO: implement a simple reset generator: it drives one reset pulse of 3cc / simulation
 
 // TODO: instantiate the ex_input_if
 // TODO: instantiate the ex_output_if
  
 // TODO: connect interfaces to clk and reset 
 // TODO: connect other wires to the interfaces
 
 // TODO: create an instance of the P2S
 // TODO: connect the instance to the clock reset and other signals
 
endmodule
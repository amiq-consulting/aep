/******************************************************************************
Copyright (c) 2004-2017, AMIQ Consulting srl. All rights reserved.

Licensed under the Apache License, Version 2.0 (the "License");
you may not use this file except in compliance with the License.
You may obtain a copy of the License at
    http://www.apache.org/licenses/LICENSE-2.0

Unless required by applicable law or agreed to in writing, software
distributed under the License is distributed on an "AS IS" BASIS,
WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
See the License for the specific language governing permissions and
limitations under the License.
 *******************************************************************************/

`ifndef __ex_out_agent
`define __ex_out_agent

/**
 * TODO: declare a class called ex_out_agent
 * Declare a field of type ex_out_monitor inside the agent which is created in the constructor
 * 
 * 
 * TODO: implement a method called set_virtual_if(virtual interface ex_in_intf aif)
 * This method must set the virtual interface fields in the driver and monitor
 * 
 */


`endif


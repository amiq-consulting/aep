/******************************************************************************
Copyright (c) 2004-2017, AMIQ Consulting srl. All rights reserved.

Licensed under the Apache License, Version 2.0 (the "License");
you may not use this file except in compliance with the License.
You may obtain a copy of the License at
    http://www.apache.org/licenses/LICENSE-2.0

Unless required by applicable law or agreed to in writing, software
distributed under the License is distributed on an "AS IS" BASIS,
WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
See the License for the specific language governing permissions and
limitations under the License.
 *******************************************************************************/
 
`ifndef __ex_scoreboard
`define __ex_scoreboard

/**
 * TODO: define the ex_scoreboard class 
 *
 * 
 * TODO: implement these tasks:
 * - listen_input() waits for new items recovered on the input interface
 * - listen_output() waits for new items recovered on the output interface  
 * 
 * TODO: implement the checking mechanism
 * 
 * TODO: implement functional coverage that target checked data
 * 
 */
 


`endif
 
